module systemTasks(input [7:0] x, output [7:0] z);
	
	assign z = ~x;

endmodule