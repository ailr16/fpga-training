module left_rotate8 (input wire clk, output wire [7:0] parallel_output);
	
endmodule 